module packet_rx(

);


endmodule
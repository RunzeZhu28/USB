module packet_tx(

);


endmodule
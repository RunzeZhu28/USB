module usb(
	output a
);

assign a =1'b1;
endmodule
module transaction(

);


endmodule